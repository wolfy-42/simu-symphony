-----------------------------------------------------------------------------
--
-- Copyright (C) 2019 Fidus Systems Inc.
--
-- Project       : RIPL 
-- Author        : Jacob von Chorus
-- Created       : 2019-02-14
-----------------------------------------------------------------------------
-----------------------------------------------------------------------------
-- Description   : Empty design unit so that xsim has a work.glbl design unit to load.
-- Updated       : date / author - comment
-----------------------------------------------------------------------------

entity glbl is
end entity glbl;

architecture rtl of glbl is
begin
end architecture rtl;
